
examples asap
