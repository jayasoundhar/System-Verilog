module str_1;
  string A="DESIGN ENGINEER";
  initial begin
    $display("A=%d",A.len);
  end
endmodule


// A= 15
