class sample;
  
  rand int a;
  rand int b[4:0];
endclass

module tb;
  sample s;
  initial begin
    s = new();
  repeat(10) begin
     s.randomize();
    $display("a=>%d\tb=>%p\t",s.a,s.b);
  end
  end
  
endmodule


a=> -384116807	b=>'{-1593209748, -1589970777, -1333235549, 2063212956, -816528844} 	
a=> 1637914715	b=>'{1233360000, 1959907722, 1981917762, 544271061, 1115228545} 	
a=>  397247290	b=>'{-277685674, 1541889331, -1282256434, 2145167130, 986512640} 	
a=> -407577593	b=>'{-1435914926, 1483337049, -1361658139, 547650128, -1635431754} 	
a=>-1298805792	b=>'{-1452694196, -907768476, -222450708, 1529991033, -2115737025} 	
a=>  842439123	b=>'{150072278, -1397549008, 1595207985, 298565361, 717502027} 	
a=> 1249691690	b=>'{1815877660, 40671725, -876975237, -2006500183, 1083171501} 	
a=> -872730637	b=>'{-354697074, -1895365839, 917123802, 449271490, -1127639830} 	
a=> 1274975648	b=>'{1343686035, 1739827842, 242394827, -586684915, 1924666731} 	
a=> 2069063609	b=>'{2014635271, -59470792, -1521330610, 1867465141, 497057233} 
