module str_1;
  string A="DESIGN ENGINEER";
  initial begin
    $display("output A=%d",A.len);
  end
endmodule


result output_str_1
KERNEL: output A= 15
