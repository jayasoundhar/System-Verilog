128123456789
