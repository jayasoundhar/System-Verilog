class sample;
  
  rand byte a;
  rand byte b[4:0];
endclass

module tb;
  sample s;
  initial begin
    s = new();
  repeat(10) begin
    s.randomize();
    $display("a=>%d\tb=>%p\t",s.a,s.b);
    s.a.rand_mode(0);
    $display("a=>%d\tb=>%p\t",s.a,s.b);
    s.randomize();
    $display("a=>%d\tb=>%p\t",s.a,s.b); 
    s.a.rand_mode(1);   
    s.randomize();
    $display("a=>%d\tb=>%p\t",s.a,s.b);
    s.randomize();
    $display("a=>%d\tb=>%p\t",s.a,s.b);
  end
  end
  
endmodule

a=>        -71	b=>'{108, -89, -93, -100, 52} 	
a=>        -71	b=>'{108, -89, -93, -100, 52} 	
a=>        -71	b=>'{91, -128, -118, 66, -43} 	
a=>         58	b=>'{86, 51, -50, 26, 0} 	
a=>          7	b=>'{82, 89, -27, 80, -74} 	
a=>        -32	b=>'{76, 100, -20, 121, 63} 	
a=>        -32	b=>'{76, 100, -20, 121, 63} 	
a=>        -32	b=>'{-45, -42, 48, 49, -15} 	
a=>         42	b=>'{28, -19, 123, -87, -83} 	
a=>        -13	b=>'{-114, 49, -38, -62, -22} 	
a=>        -96	b=>'{-109, -126, -53, 13, 107} 	
a=>        -96	b=>'{-109, -126, -53, 13, 107} 	
a=>        -96	b=>'{-71, 7, 56, 78, -75} 	
a=>        -75	b=>'{-85, -90, 56, -4, -9} 	
a=>        -16	b=>'{66, -1, -60, 7, -78} 	
a=>         99	b=>'{3, 12, 6, -29, 54} 	
a=>         99	b=>'{3, 12, 6, -29, 54} 	
a=>         99	b=>'{26, 14, -99, -79, -23} 	
a=>        -11	b=>'{-124, -1, -20, -55, 34} 	
a=>       -102	b=>'{-16, 12, -110, -50, 42} 	
a=>        -90	b=>'{35, -105, 26, -52, 15} 	
a=>        -90	b=>'{35, -105, 26, -52, 15} 	
a=>        -90	b=>'{0, -85, -49, -69, -98} 	
a=>        -31	b=>'{98, -53, -29, -115, 73} 	
a=>          6	b=>'{-59, -67, 7, -70, 36} 	
a=>         47	b=>'{-95, 58, -6, 78, -22} 	
a=>         47	b=>'{-95, 58, -6, 78, -22} 	
a=>         47	b=>'{-125, -44, 100, 33, -62} 	
a=>        116	b=>'{-25, -21, -31, 116, -13} 	
a=>       -112	b=>'{-105, 86, -126, 80, 87} 	
a=>         91	b=>'{-101, -116, -27, -40, 73} 	
a=>         91	b=>'{-101, -116, -27, -40, 73} 	
a=>         91	b=>'{-32, -123, 20, 116, -57} 	
a=>        -24	b=>'{-74, 67, -83, -4, 111} 	
a=>         33	b=>'{-93, 84, 40, 123, -63} 	
a=>        -78	b=>'{-53, -13, -74, 0, -49} 	
a=>        -78	b=>'{-53, -13, -74, 0, -49} 	
a=>        -78	b=>'{-105, -3, -127, -107, 82} 	
a=>        -53	b=>'{125, -38, -30, -98, 111} 	
a=>         78	b=>'{-114, 119, 78, -96, 0} 	
a=>        109	b=>'{-93, 56, -119, 23, -126} 	
a=>        109	b=>'{-93, 56, -119, 23, -126} 	
a=>        109	b=>'{-52, -11, -38, -110, -56} 	
a=>          9	b=>'{-58, 10, 47, 78, -53} 	
a=>         81	b=>'{0, 116, -13, 73, 63} 	
a=>        -20	b=>'{-88, 68, 10, -10, -95} 	
a=>        -20	b=>'{-88, 68, 10, -10, -95} 	
a=>        -20	b=>'{68, -30, 20, -98, 1} 	
a=>        -14	b=>'{-124, -45, 127, -12, -41} 	
a=>         96	b=>'{-26, -98, 115, 54, -3} 
