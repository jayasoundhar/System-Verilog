module str_02;
  string A =("design_engineer");
  initial begin
  $display("yours output on A=%s ",A.toupper());
  end
endmodule

results
KERNEL: yours output's str_02 on A=DESIGN_ENGINEER
