module str_05;
  string A=("DESIGN_ENGINEER");
  initial begin
    $display("A=%s",A.getc(2));
  end
endmodule

// E
