module str_06;
  string A=("3455647RING");
  initial begin
    $display("A=%d",A.atoi());
  end
endmodule

// 3455647
