module str_06;
  string A=("3455647RING");
  initial begin
    $display("your's expected output for str_06 is A=%d",A.atoi());
  end
endmodule

result
KERNEL: your's expected output for str_06 is A=    3455647
