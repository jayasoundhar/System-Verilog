123456778990
