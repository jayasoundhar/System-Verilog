
module str_11;
  string A="DESIGN";
  initial begin
    $display("A =%s",A.substr(2,3));
  end
endmodule


// A =SI
