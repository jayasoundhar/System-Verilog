module str_02;
  string A =("design_engineer");
  initial begin
  $display("A=%s ",A.toupper());
  end
endmodule

// A=DESIGN_ENGINEER
